`timescale 1ns / 1ps

module uart #(
    parameter LOGD = 7
  ) (
    input wire                     clk,
    input wire                     i_reset,
    input wire                     wr_valid,
    // verilator lint_off UNUSEDSIGNAL
    input wire  [31:0]             wr_data,
    // verilator lint_on UNUSEDSIGNAL
    input wire  [31:0]             wr_addr,
    output wire                    uart_rxd_out
  );

  wire   tx_valid;
  assign tx_valid = wr_valid && wr_addr[LOGD];

  tx txi (
    clk,
    i_reset,
    tx_valid,
    wr_data[7:0],
    uart_rxd_out
  );
endmodule
